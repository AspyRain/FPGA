
`ifndef DEFINES_VH
`define DEFINES_VH
`define T0H 4'd15
`define T0L 4'd40
`define T1H 4'd40
`define T1L 4'd40
`define RST 14'd15_000
//GRB 24bit ，高位先发(msb)
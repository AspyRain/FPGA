module counter_key (
    input           clk     ,
    input           rst_n   ,
    output [16:0]   dout    ,
    input           key     ,
    output     reg      flag    
);





endmodule

